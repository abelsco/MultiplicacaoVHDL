library verilog;
use verilog.vl_types.all;
entity CODE8B_vlg_vec_tst is
end CODE8B_vlg_vec_tst;
